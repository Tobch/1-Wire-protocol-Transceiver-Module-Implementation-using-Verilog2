`timescale 1ns/1ps

//------------------------------------------------------------------------------
// File: one_wire_timing.v
//------------------------------------------------------------------------------
module one_wire_timing (
    input clk,
    input rst_n
);
    // purely parameter container
endmodule