`timescale 1ns/1ps

//------------------------------------------------------------------------------
// File: one_wire_timing.v
// Description: Parameter definitions for 1-Wire protocol timing (standard speed)
//------------------------------------------------------------------------------
module one_wire_timing (
    input clk,
    input rst_n
);
    // purely parameter container
endmodule